`timescale 1ns / 1ps

module ExceptionUnit (
    input clk,
    rst,
    input csr_rw_in,
    // write/set/clear (funct bits from instruction)
    input [1:0] csr_wsc_mode_in,
    input csr_w_imm_mux,
    input [11:0] csr_rw_addr_in,
    input [31:0] csr_w_data_reg,
    input [4:0] csr_w_data_imm,
    output [31:0] csr_r_data_out,

    input interrupt,
    input illegal_inst,
    input l_access_fault,
    input s_access_fault,
    input ecall_m,

    input mret,

    input [31:0] epc_cur,
    input [31:0] epc_next,
    output [31:0] PC_redirect,
    output redirect_mux,

    output reg_FD_flush,
    reg_DE_flush,
    reg_EM_flush,
    reg_MW_flush,
    output RegWrite_cancel,
    output MemWrite_cancel
);
  // According to the diagram, design the Exception Unit
  // You can modify any code in this file if needed!
  reg [11:0] csr_waddr;
  reg [31:0] csr_wdata;
  reg csr_w;
  reg [1:0] csr_wsc;
  wire [11:0] csr_raddr;

  wire [31:0] mstatus;
  wire [31:0] csr_rdata;

  CSRRegs csr (
      .clk(clk),
      .rst(rst),
      .csr_w(csr_w),
      .raddr(csr_raddr),
      .waddr(csr_waddr),
      .wdata(csr_wdata),
      .rdata(csr_rdata),
      .mstatus(mstatus),
      .csr_wsc_mode(csr_wsc)
  );



endmodule
